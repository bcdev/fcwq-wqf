netcdf in {
dimensions:
	time = 8 ;
	lat = 469 ;
	lon = 527 ;
variables:
	float chl(time, lat, lon) ;
		chl:_FillValue = NaNf ;
		string chl:standard_name = "chlorophyll_concentration_in_sea_water" ;
		string chl:units = "mg m-3" ;
		chl:_Storage = "chunked" ;
		chl:_ChunkSizes = 8, 67, 31 ;
		chl:_DeflateLevel = 1 ;
		chl:_Shuffle = "true" ;
		chl:_Endianness = "little" ;
	float deptho(lat, lon) ;
		deptho:_FillValue = NaNf ;
		string deptho:standard_name = "sea_floor_depth_below_geoid" ;
		string deptho:units = "m" ;
		deptho:_Storage = "chunked" ;
		deptho:_ChunkSizes = 67, 31 ;
		deptho:_DeflateLevel = 1 ;
		deptho:_Shuffle = "true" ;
		deptho:_Endianness = "little" ;
	float doy(time) ;
		doy:_FillValue = NaNf ;
		string doy:long_name = "day of year" ;
		doy:_Storage = "contiguous" ;
		doy:_Endianness = "little" ;
	float mdt(lat, lon) ;
		mdt:_FillValue = NaNf ;
		string mdt:standard_name = "sea_surface_height_above_geoid" ;
		string mdt:units = "m" ;
		mdt:_Storage = "chunked" ;
		mdt:_ChunkSizes = 67, 31 ;
		mdt:_DeflateLevel = 1 ;
		mdt:_Shuffle = "true" ;
		mdt:_Endianness = "little" ;
	float mlotst(time, lat, lon) ;
		mlotst:_FillValue = NaNf ;
		string mlotst:standard_name = "ocean_mixed_layer_thickness_defined_by_sigma_theta" ;
		string mlotst:units = "m" ;
		mlotst:_Storage = "chunked" ;
		mlotst:_ChunkSizes = 8, 67, 31 ;
		mlotst:_DeflateLevel = 1 ;
		mlotst:_Shuffle = "true" ;
		mlotst:_Endianness = "little" ;
	float no3(time, lat, lon) ;
		no3:_FillValue = NaNf ;
		string no3:standard_name = "mole_concentration_of_nitrate_in_sea_water" ;
		string no3:units = "mmol m-3" ;
		no3:_Storage = "chunked" ;
		no3:_ChunkSizes = 8, 67, 31 ;
		no3:_DeflateLevel = 1 ;
		no3:_Shuffle = "true" ;
		no3:_Endianness = "little" ;
	float o2(time, lat, lon) ;
		o2:_FillValue = NaNf ;
		string o2:standard_name = "mole_concentration_of_dissolved_molecular_oxygen_in_sea_water" ;
		string o2:units = "mmol m-3" ;
		o2:_Storage = "chunked" ;
		o2:_ChunkSizes = 8, 67, 31 ;
		o2:_DeflateLevel = 1 ;
		o2:_Shuffle = "true" ;
		o2:_Endianness = "little" ;
	float ph(time, lat, lon) ;
		ph:_FillValue = NaNf ;
		string ph:standard_name = "sea_water_ph_reported_on_total_scale" ;
		string ph:units = "1" ;
		ph:_Storage = "chunked" ;
		ph:_ChunkSizes = 8, 67, 31 ;
		ph:_DeflateLevel = 1 ;
		ph:_Shuffle = "true" ;
		ph:_Endianness = "little" ;
	float po4(time, lat, lon) ;
		po4:_FillValue = NaNf ;
		string po4:standard_name = "mole_concentration_of_phosphate_in_sea_water" ;
		string po4:units = "mmol m-3" ;
		po4:_Storage = "chunked" ;
		po4:_ChunkSizes = 8, 67, 31 ;
		po4:_DeflateLevel = 1 ;
		po4:_Shuffle = "true" ;
		po4:_Endianness = "little" ;
	float so(time, lat, lon) ;
		so:_FillValue = NaNf ;
		string so:standard_name = "sea_water_salinity" ;
		string so:units = "1e-3" ;
		so:_Storage = "chunked" ;
		so:_ChunkSizes = 8, 67, 31 ;
		so:_DeflateLevel = 1 ;
		so:_Shuffle = "true" ;
		so:_Endianness = "little" ;
	float ssrd(time, lat, lon) ;
		ssrd:_FillValue = NaNf ;
		string ssrd:standard_name = "surface_downwelling_shortwave_flux_in_air" ;
		string ssrd:units = "J m**-2" ;
		ssrd:_Storage = "chunked" ;
		ssrd:_ChunkSizes = 8, 67, 31 ;
		ssrd:_DeflateLevel = 1 ;
		ssrd:_Shuffle = "true" ;
		ssrd:_Endianness = "little" ;
	float sst(time, lat, lon) ;
		sst:_FillValue = NaNf ;
		string sst:long_name = "Sea surface temperature" ;
		string sst:units = "K" ;
		sst:_Storage = "chunked" ;
		sst:_ChunkSizes = 8, 67, 31 ;
		sst:_DeflateLevel = 1 ;
		sst:_Shuffle = "true" ;
		sst:_Endianness = "little" ;
	float tcc(time, lat, lon) ;
		tcc:_FillValue = NaNf ;
		string tcc:standard_name = "cloud_area_fraction" ;
		string tcc:units = "(0 - 1)" ;
		tcc:_Storage = "chunked" ;
		tcc:_ChunkSizes = 8, 67, 31 ;
		tcc:_DeflateLevel = 1 ;
		tcc:_Shuffle = "true" ;
		tcc:_Endianness = "little" ;
	float thetao(time, lat, lon) ;
        thetao:_FillValue = NaNf ;
        string thetao:long_name = "Sea Water Potential Temperature" ;
        string thetao:standard_name = "sea_water_potential_temperature" ;
        string thetao:units = "degrees_C" ;
        thetao:_Storage = "chunked" ;
        thetao:_ChunkSizes = 8, 67, 31 ;
        thetao:_Shuffle = "true" ;
        thetao:_DeflateLevel = 1 ;
        thetao:_Endianness = "little" ;
	float tp(time, lat, lon) ;
		tp:_FillValue = NaNf ;
		string tp:long_name = "Total precipitation" ;
		string tp:units = "m" ;
		tp:_Storage = "chunked" ;
		tp:_ChunkSizes = 8, 67, 31 ;
		tp:_DeflateLevel = 1 ;
		tp:_Shuffle = "true" ;
		tp:_Endianness = "little" ;
	float u10(time, lat, lon) ;
		u10:_FillValue = NaNf ;
		string u10:long_name = "10 metre U wind component" ;
		string u10:units = "m s**-1" ;
		u10:_Storage = "chunked" ;
		u10:_ChunkSizes = 8, 67, 31 ;
		u10:_DeflateLevel = 1 ;
		u10:_Shuffle = "true" ;
		u10:_Endianness = "little" ;
	float uo(time, lat, lon) ;
		uo:_FillValue = NaNf ;
		string uo:standard_name = "eastward_sea_water_velocity" ;
		string uo:units = "m s-1" ;
		uo:_Storage = "chunked" ;
		uo:_ChunkSizes = 8, 67, 31 ;
		uo:_DeflateLevel = 1 ;
		uo:_Shuffle = "true" ;
		uo:_Endianness = "little" ;
	float v10(time, lat, lon) ;
		v10:_FillValue = NaNf ;
		string v10:long_name = "10 metre V wind component" ;
		string v10:units = "m s**-1" ;
		v10:_Storage = "chunked" ;
		v10:_ChunkSizes = 8, 67, 31 ;
		v10:_DeflateLevel = 1 ;
		v10:_Shuffle = "true" ;
		v10:_Endianness = "little" ;
	float vo(time, lat, lon) ;
		vo:_FillValue = NaNf ;
		string vo:standard_name = "northward_sea_water_velocity" ;
		string vo:units = "m s-1" ;
		vo:_Storage = "chunked" ;
		vo:_ChunkSizes = 8, 67, 31 ;
		vo:_DeflateLevel = 1 ;
		vo:_Shuffle = "true" ;
		vo:_Endianness = "little" ;
	float zos(time, lat, lon) ;
		zos:_FillValue = NaNf ;
		string zos:standard_name = "sea_surface_height_above_geoid" ;
		string zos:units = "m" ;
		zos:_Storage = "chunked" ;
		zos:_ChunkSizes = 8, 67, 31 ;
		zos:_DeflateLevel = 1 ;
		zos:_Shuffle = "true" ;
		zos:_Endianness = "little" ;
	double lat(lat) ;
		lat:_FillValue = NaN ;
		string lat:standard_name = "latitude" ;
		string lat:units = "degrees_north" ;
		lat:_Storage = "contiguous" ;
		lat:_Endianness = "little" ;
	double lon(lon) ;
		lon:_FillValue = NaN ;
		string lon:standard_name = "longitude" ;
		string lon:units = "degrees_east" ;
		lon:_Storage = "contiguous" ;
		lon:_Endianness = "little" ;
	double time(time) ;
		time:_FillValue = NaN ;
		string time:_CoordinateAxisType = "Time" ;
		string time:axis = "T" ;
		string time:standard_name = "time" ;
		string time:units = "days since 2020-07-01 00:00:00" ;
		string time:calendar = "proleptic_gregorian" ;
		time:_Storage = "contiguous" ;
		time:_Endianness = "little" ;

// global attributes:
		:_NCProperties = "version=2,h5netcdf=1.3.0,hdf5=1.14.3,h5py=3.11.0" ;
		:_SuperblockVersion = 0 ;
		:_IsNetcdf4 = 1 ;
		:_Format = "netCDF-4" ;
}
